module 



endmodule