
module testbench();

	reg 
	wire 
	
	//Ejercicio #1
	
	tabla_1 T1(p1,p2,p3,p4,led1);
	
	tabla_2 T2(p4,led2);
	
	tabla_3 T3(p5,p6,p7,p8,led3);
	
	tabla_4 T4(p9,p10,p11,p12,led4);
	
	//	Ejercicio #2 
	
	tabla_1_2 T1_2(p13,p14,p15,p16,led5);
	
	tabla_2_2 T2_2(p17,p18,led6);
	
	tabla_3_2 T3_2(p19,p20,led7);
	
	tabla_4_2 T4_2(p21,p22,led8);
	
	initial begin
		
		$display();